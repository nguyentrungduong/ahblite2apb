////////////////////////////////////////////////////////////////////////////////
// Company     : SH Consulting
//
// Filename    : mux16.v
// Description : 16:1 parallel mux.
//
// Author      : Duong Nguyen
// Created On  : 10-6-2015
// History     : Initial 	
//
////////////////////////////////////////////////////////////////////////////////

module mux16
    (
    sel0,
    in0,
    //-------------------
    sel1,
    in1,
    //-------------------
    sel2,
    in2,
    //-------------------
    sel3,
    in3,
    //-------------------
    sel4,
    in4,
    //-------------------
    sel5,
    in5,
    //-------------------
    sel6,
    in6,
    //-------------------
    sel7,
    in7,
    //-------------------
    sel8,
    in8,
    //-------------------
    sel9,
    in9,
    //-------------------
    sel10,
    in10,
    //-------------------
    sel11,
    in11,
    //-------------------
    sel12,
    in12,
    //-------------------
    sel13,
    in13,
    //-------------------
    sel14,
    in14,
    //-------------------
    sel15,
    in15,
    //-------------------
    out
    );

//------------------------------------------------------------------------------
//Parameters
parameter DW = 1'b1;
//------------------------------------------------------------------------------
// Port declarations
input               sel0;
input [DW-1:0]	    in0;
//
input               sel1;
input [DW-1:0]	    in1;
//
input               sel2;
input [DW-1:0]	    in2;
//
input               sel3;
input [DW-1:0]	    in3;
//
input               sel4;
input [DW-1:0]	    in4;
//
input               sel5;
input [DW-1:0]	    in5;
//
input               sel6;
input [DW-1:0]	    in6;
//
input               sel7;
input [DW-1:0]	    in7;
//
input               sel8;
input [DW-1:0]	    in8;
//
input               sel9;
input [DW-1:0]	    in9;
//
input               sel10;
input [DW-1:0]	    in10;
//
input               sel11;
input [DW-1:0]	    in11;
//
input               sel12;
input [DW-1:0]	    in12;
//
input               sel13;
input [DW-1:0]	    in13;
//
input               sel14;
input [DW-1:0]	    in14;
//
input               sel15;
input [DW-1:0]	    in15;
//
output [DW-1:0]	    out;
//------------------------------------------------------------------------------
//internal signal
wire [DW-1:0]       out0_7;
wire [DW-1:0]       out8_15;
//------------------------------------------------------------------------------
//Mux 8:1
mux8   #(.DW(DW))   mux0_7
    (
    .sel0  (sel0),
    .in0   (in0),
    //-------------------
    .sel1  (sel1),
    .in1   (in1),
    //-------------------
    .sel2  (sel2),
    .in2   (in2),
    //-------------------
    .sel3  (sel3),
    .in3   (in3),
    //-------------------
    .sel4  (sel4),
    .in4   (in4),
    //-------------------
    .sel5  (sel5),
    .in5   (in5),
    //-------------------
    .sel6  (sel6),
    .in6   (in6),
    //-------------------
    .sel7  (sel7),
    .in7   (in7),
    //-------------------
    .out   (out0_7)
    );
//------------------------------------------------------------------------------
//Mux 8:1
mux8   #(.DW(DW))   mux8_15
    (
    .sel0  (sel8),
    .in0   (in8),
    //-------------------
    .sel1  (sel9),
    .in1   (in9),
    //-------------------
    .sel2  (sel10),
    .in2   (in10),
    //-------------------
    .sel3  (sel11),
    .in3   (in11),
    //-------------------
    .sel4  (sel12),
    .in4   (in12),
    //-------------------
    .sel5  (sel13),
    .in5   (in13),
    //-------------------
    .sel6  (sel14),
    .in6   (in14),
    //-------------------
    .sel7  (sel15),
    .in7   (in15),
    //-------------------
    .out   (out8_15)
    );
//------------------------------------------------------------------------------
//Mux 2:1
assign out = out0_7 | out8_15;

endmodule 

